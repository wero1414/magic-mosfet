magic
tech sky130A
timestamp 1612038143
<< nmos >>
rect 40 0 55 65
<< ndiff >>
rect 0 45 40 65
rect 0 25 6 45
rect 25 25 40 45
rect 0 0 40 25
rect 55 40 95 65
rect 55 15 70 40
rect 90 15 95 40
rect 55 0 95 15
<< ndiffc >>
rect 6 25 25 45
rect 70 15 90 40
<< poly >>
rect 40 65 55 110
rect 40 -20 55 0
rect -5 -30 55 -20
rect -5 -49 10 -30
rect 30 -49 55 -30
rect -5 -55 55 -49
<< polycont >>
rect 10 -49 30 -30
<< locali >>
rect -54 45 30 65
rect -54 25 -50 45
rect -25 25 6 45
rect 25 25 30 45
rect -54 0 30 25
rect 65 40 155 50
rect 65 15 70 40
rect 90 38 155 40
rect 90 21 130 38
rect 150 21 155 38
rect 90 15 155 21
rect 65 4 155 15
rect -50 -30 35 -20
rect -50 -50 -45 -30
rect -24 -49 10 -30
rect 30 -49 35 -30
rect -24 -50 35 -49
rect -50 -60 35 -50
<< viali >>
rect -50 25 -25 45
rect 130 21 150 38
rect -45 -50 -24 -30
<< metal1 >>
rect -145 45 -15 50
rect -145 25 -50 45
rect -25 25 -15 45
rect -145 20 -15 25
rect 125 38 220 45
rect 125 21 130 38
rect 150 21 220 38
rect 125 15 220 21
rect -120 -30 -15 -25
rect -120 -50 -45 -30
rect -24 -50 -15 -30
rect -120 -55 -15 -50
rect -119 -56 -15 -55
<< labels >>
rlabel metal1 -140 25 -121 45 1 source
rlabel metal1 -115 -49 -90 -30 1 gate
rlabel metal1 190 20 215 40 1 drain
<< end >>
